`timescale 1ns / 1ps
`include "../../incl.vh"

//
// Memory instances of XPHM
//
module xphm_mem (
    input clk,
    // Read ports
    input rd_en,
    input [$clog2(`XPHM_DEPTH)-1:0] rd_addr,
    output [`XPHM_DATA_WIDTH-1:0] dout,
    // Write ports
    input wr_en,
    input [$clog2(`XPHM_DEPTH)-1:0] wr_addr,
    input [`XPHM_DATA_WIDTH-1:0] din
);
    sdp_bram #(
        .DATA_WIDTH(`XPHM_DATA_WIDTH),
        .DEPTH(`XPHM_DEPTH),
        .NUM_PIPE(`XPHM_NUM_PIPE)
    ) sdp_bram_inst(
    	.clk(clk),
        .wr_en(wr_en),
        .din(din),
        .wr_addr(wr_addr),
        .rd_en(rd_en),
        .rd_addr(rd_addr),
        .dout(dout)
    );
endmodule
