//
// This file is a configuration file.
// It can not be included directly. 
// We should use tools/gen_incl.py to generate a new verilog header file which can be included.
//

// Hyper Parameters
`define M 32
`define P 96
`define Q 16
`define R 16
`define S 8

// `define DEBUG

// Instruction type definition
`define INS_NONE 8'b11111111
`define INS_CONV 8'b00000001
`define INS_MAXP 8'b00000010
`define INS_AVGP 8'b00000011
`define INS_ADD 8'b00000100
`define INS_REMAP 8'b00000101
`define INS_FC 8'b00000110

// RTM (URAM)
// Data width: S*R*8
`define RTM_DEPTH 65536
`define RTM_URAM_NUM_PIPE 11

// CWM (URAM)
// Data width: M*4*8
`define CWM_DEPTH 163840
`define CWM_NUM_PIPE 14

// IM (BRAM)
`define INS_RAM_DATA_WIDTH 512
`define INS_RAM_DEPTH 1024
`define INS_RAM_NUM_PIPE 3

// BM (BRAM)
`define BM_DATA_WIDTH 512
`define BM_DEPTH 8192
`define BM_NUM_PIPE 2

// XPHM (BRAM)
`define XPHM_X_a__WIDTH 16
`define XPHM_len_per_chan_WIDTH 16
`define XPHM_win_x_WIDTH 16
`define XPHM_win_y_WIDTH 16
`define XPHM_DATA_WIDTH (`XPHM_X_a__WIDTH+`XPHM_len_per_chan_WIDTH+`XPHM_win_x_WIDTH+`XPHM_win_y_WIDTH)
`define XPHM_DEPTH 8192
`define XPHM_NUM_PIPE 2

// MXM (URAM)
// Data width: P*2*8
`define MXM_DEPTH 8192
`define MXM_PROG_FULL (`MXM_DEPTH-32)
`define MXM_NUM_PIPE 4

// X-bus
`define XBUS_TAG_WIDTH 2
`define XBUS_TAG_INVALID 0
`define XBUS_TAG_HEAD 1
`define XBUS_TAG_BODY 2
`define XBUS_TAG_END 3
`define XBUS_CACHE_DEPTH 512
`define XBUS_CACHE_FULL 256

// Systolic Array
`define SA_TAG_DW 1
`define SA_TAG_END 1'b1
`define SA_TAG_NONE 1'b0

`define LATENCY_COUNTER_WIDTH 32

// XDMA
`define XDMA_USR_INTR_COUNT 16
`define XDMA_AXIS_DATA_WIDTH 512
`define XDMA_AXIS_KEEP_WIDTH (`XDMA_AXIS_DATA_WIDTH/8)

// sr_cr AXI4LITE
`define SR_CR_AXI_ADDR_WIDTH 8
`define SR_CR_AXI_DATA_WIDTH 32

// DMA AXI IF
`define DMA_AXI_DATA_WIDTH 512
`define DDR_AXI_ADDR_WIDTH 32
`define DDR_AXI_STRB_WIDTH 64
`define DDR_AXI_ID_WIDTH 8
`define DDR_AXI_MAX_BURST_LEN 256
`define DDR_AXIS_DATA_WIDTH 512
`define DDR_AXIS_KEEP_ENABLE 1
`define DDR_AXIS_KEEP_WIDTH 64
`define DDR_AXIS_LAST_ENABLE 1
`define DDR_AXIS_ID_ENABLE 0
`define DDR_AXIS_ID_WIDTH 8
`define DDR_AXIS_DEST_ENABLE 0
`define DDR_AXIS_DEST_WIDTH 8
`define DDR_AXIS_USER_ENABLE 0
`define DDR_AXIS_USER_WIDTH 1
`define DDR_LEN_WIDTH 27
`define DDR_TAG_WIDTH 8
